LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY LZE IS
PORT( LZE_IN   : in STD_LOGIC_VECTOR(31 DOWNTO 0);
		LZE_OUT  : out STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END ENTITY;

ARCHITECTURE Behavior OF LZE IS
SIGNAL zeros: STD_LOGIC_VECTOR(15 DOWNTO 0) := (others => '0');
BEGIN
	LZE_out <= zeros & LZE_in(15 DOWNTO 0);
END Behavior;

